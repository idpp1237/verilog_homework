module InstructionMemory(
Addr_in,
instr);
input [31:0]Addr_in;
output reg[31:0]instr; 

always@(*)
begin
case(Addr_in)

0:instr=32'b010100_01100_01101_01011_00000_011011;//
4:instr=32'b010100_01001_01010_01000_00000_001001;//
8:instr=32'b010100_01001_01010_01001_00000_010010;//
12:instr=32'b000000_00000_00000_00000_00000_000000;	//stall			//stall
16:instr=32'b010100_01011_01111_01101_00000_100100;//

20:instr=32'b101001_01011_01000_00000_00000_000010;
24:instr=32'b101010_01011_10011_00000_00000_000010;
//
28:instr=32'b101001_01010_10100_00000_00000_000100;
32:instr=32'b101001_01010_01000_00000_00000_000010;
36:instr=32'b101010_01011_10100_00000_00000_000011;
40:instr=32'b101000_10000_10111_00000_00000_000010;
44:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
48:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
52:instr=32'b100111_10100_10101_00000_00000_101000;
56:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
60:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
64:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
68:instr=32'b100111_10101_10110_00000_00000_010110; 
72:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
76:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
80:instr=32'b000000_00000_00000_00000_00000_000000;	//stall
84:instr=32'b101000_10110_10011_00000_00000_001000; 
							




default :instr=32'b0;
endcase
end
endmodule
