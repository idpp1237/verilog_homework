module InstructionMemory(
Addr_in,
instr);
input [31:0]Addr_in;
output reg[31:0]instr; 

always@(*)
begin
case(Addr_in)
0:instr=32'b0101_0001_0010_1010_0100_0000_0000_1001;
4:instr=32'b0101_0001_0010_1010_0100_1000_0001_0010;
8:instr=32'b0101_0001_1000_1101_0101_1000_0001_1011;
12:instr=32'b0101_0001_1100_1111_0110_1000_0010_0100;
16:instr=32'b1010_0101_0110_1000_0000_0000_0000_0010;
20:instr=32'b10101001011100110000000000000010;
24:instr=32'b10101001011101000000000000000011;
28:instr=32'b10100101010010000000000000000010;
32:instr=32'b10100101010101000000000000000100;
36:instr=32'b10011110100101010000000000101000;
40:instr=32'b10011110101101100000000000010110; 
44:instr=32'b10100010110100110000000000001000; 
48:instr=32'b10100010000101110000000000000010;
52:instr=32'b01110001110011000000000000000100;
56:instr=32'b01110011000011000000000000000100;
60:instr=32'b01110010101100110000000000000100;
64:instr=32'b01110011001110000000000000000100;
68:instr=32'b01101100000000000000000001101110;
default :instr=32'b0;
endcase
end
endmodule
